`timescale 1ns / 1ps
`include "../src/mips/mips_pkg.vh"

module mips_simple_tb();

  // Señales para conectar al DUT
  reg clk;
  reg reset;
  wire [`DATA_WIDTH-1:0] result;
  wire halt;  // Agregamos un wire para la señal de halt
  
  // Instancia del módulo MIPS
  mips dut (
    .clk    (clk),
    .reset  (reset),
    .result (result),
    .halt   (halt),  // Conectamos la señal de halt para detectar fin de ejecución
    .stall  (1'b0)   // No se usa stall en este testbench
  );
  
  // Genera un reloj de 10ns (100 MHz)
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end
  
  // Variables para el ciclo
  integer cycle_count;
  
  // Función para mostrar el tipo de instrucción
  function [8*20:1] instr_type;
    input [`DATA_WIDTH-1:0] instr;
    reg [5:0] opcode;
    begin
      opcode = instr[31:26];
      case(opcode)
        `OPCODE_R_TYPE: instr_type = "R-type";
        `OPCODE_ADDI:   instr_type = "addi";
        `OPCODE_LW:     instr_type = "lw";
        `OPCODE_SW:     instr_type = "sw";
        `OPCODE_BEQ:    instr_type = "beq";
        `OPCODE_BNE:    instr_type = "bne";
        default:        instr_type = "desconocida";
      endcase
    end
  endfunction
  
  // Inicio de la simulación
  initial begin
    // Inicialización de señales
    reset = 1;
    cycle_count = 0;
    
    // Mostrar encabezado
    $display("\n==== MIPS Pipeline Simple Testbench con Forwarding Unit ====\n");
    $display("Este testbench evalúa el funcionamiento del pipeline MIPS");
    $display("La simulación terminará automáticamente cuando la señal halt se active");
    
    // Liberar el reset después de unos ciclos
    #15;
    reset = 0;
    
    // Esperar hasta que halt sea 1 o hasta un tiempo máximo por seguridad
    fork
      // Opción 1: Terminar cuando halt sea 1
      begin
        wait(halt);
        $display("\n==== Procesador terminado: señal halt detectada (t=%0t ns) ====", $time);
        
        // Realizar la verificación final al detectar halt
        $display("\n==== VERIFICACIÓN FINAL AL DETECTAR HALT (Ciclo %0d) ====", cycle_count);
        $display("Registros finales:");
        $display("$1=%0d (Esperado: 5)", 
               dut.id_stage_inst.reg_bank.registers[1]);
        $display("$2=%0d (Esperado: 10)", 
               dut.id_stage_inst.reg_bank.registers[2]);
        $display("$3=%0d (Esperado: 100)", 
               dut.id_stage_inst.reg_bank.registers[3]);
        $display("$4=%0d (Esperado: 20)", 
               dut.id_stage_inst.reg_bank.registers[4]);
        $display("$5=%0d (Esperado: 5)", 
               dut.id_stage_inst.reg_bank.registers[5]);
        $display("$6=%0d (Esperado: 5)", 
               dut.id_stage_inst.reg_bank.registers[6]);
        $display("$7=%0d (Esperado: 10)", 
               dut.id_stage_inst.reg_bank.registers[7]);
        $display("$8=%0d (Esperado: 39)", 
               dut.id_stage_inst.reg_bank.registers[8]);
        $display("$9=%0d (Esperado: 1)", 
               dut.id_stage_inst.reg_bank.registers[9]);
        $display("$10=%0d", dut.id_stage_inst.reg_bank.registers[10]);
        $display("$11=%0d (Esperado: 5)", 
               dut.id_stage_inst.reg_bank.registers[11]);
        $display("$12=%0d (Esperado: 10)", 
               dut.id_stage_inst.reg_bank.registers[12]);
        $display("$13=%0d (Esperado: 0)", 
               dut.id_stage_inst.reg_bank.registers[13]);
        $display("$14=%0d (Esperado: 7)", 
               dut.id_stage_inst.reg_bank.registers[14]);
        $display("$15=%0d (Esperado: 20)", 
               dut.id_stage_inst.reg_bank.registers[15]);
               
        // Verificar memoria
        $display("\nMemoria final:");
        $display("Mem[100]=%0d (Esperado: 5)", 
               dut.mem_stage_inst.data_mem.memory[25]);
        $display("Mem[104]=%0d (Esperado: 5)", 
               dut.mem_stage_inst.data_mem.memory[26]);
        $display("Mem[35]=%0d (Esperado: 15)", 
               dut.mem_stage_inst.data_mem.memory[8]);
        $display("Mem[39]=%0d (Esperado: 35)", 
               dut.mem_stage_inst.data_mem.memory[9]);
               
        // Verificar resultado
        if (dut.id_stage_inst.reg_bank.registers[1] == 5 &&
            dut.id_stage_inst.reg_bank.registers[2] == 10 &&
            dut.id_stage_inst.reg_bank.registers[3] == 100 &&
            dut.id_stage_inst.reg_bank.registers[4] == 20 &&
            dut.id_stage_inst.reg_bank.registers[5] == 5 &&
            dut.id_stage_inst.reg_bank.registers[6] == 5 &&
            dut.id_stage_inst.reg_bank.registers[7] == 10 &&
            dut.id_stage_inst.reg_bank.registers[8] == 39 &&
            dut.id_stage_inst.reg_bank.registers[9] == 1 &&
            dut.id_stage_inst.reg_bank.registers[11] == 5 &&
            dut.id_stage_inst.reg_bank.registers[12] == 10 &&
            dut.id_stage_inst.reg_bank.registers[13] == 0 &&
            dut.id_stage_inst.reg_bank.registers[14] == 7 &&
            dut.id_stage_inst.reg_bank.registers[15] == 20 &&
            dut.mem_stage_inst.data_mem.memory[25] == 5 &&
            dut.mem_stage_inst.data_mem.memory[26] == 5 &&
            dut.mem_stage_inst.data_mem.memory[8] == 15 &&
            dut.mem_stage_inst.data_mem.memory[9] == 35) begin
          $display("\n¡PRUEBA EXITOSA! Todos los resultados son correctos.");
          $display("\nLa unidad de forwarding ha manejado correctamente los riesgos de datos resolubles.");
          $display("Los NOPs insertados han ayudado a evitar los riesgos no resolubles mediante forwarding.");
          $display("(Principalmente: load-use hazards y dependencias EX-EX que requieren stalls)");
        end else begin
          $display("\n¡PRUEBA FALLIDA! Algunos resultados no coinciden con los valores esperados.");
        end
        
        $finish;
      end
      
      // Opción 2: Tiempo máximo de seguridad
      begin
        #2000;  // Tiempo máximo de seguridad (2000 ns)
        $display("\n==== ADVERTENCIA: Se alcanzó tiempo máximo sin detectar señal halt ====");
        $finish;
      end
    join
  end
  
  // Imprime el estado de cada etapa en cada ciclo
  always @(posedge clk) begin
    if (!reset) begin
      cycle_count = cycle_count + 1;
      
      // Mostrar información del ciclo
      $display("\n==== Ciclo %0d (t=%0t ns) ====", cycle_count, $time);
      
      // Mostrar el estado del pipeline
      $display("IF: PC=%0h, Instr=%0h, Tipo=%s", 
               dut.if_stage_inst.pc_inst.pc,
               dut.if_instr,
               instr_type(dut.if_instr));
      
        $display("ID: Instr=%0h, RegDst=%0b, OpCode=%0b, ALUSrcA=%0b, ALUSrcB=%0b, Shamt=0x%h, Function=%0b, RegWrite=%0b", 
                 dut.id_instr,
                 dut.id_reg_dst,
                 dut.id_opcode,
                 dut.id_alu_src_a,
                 dut.id_alu_src_b,
                 dut.id_shamt,
                 dut.id_function,
                 dut.id_reg_write);

        $display("Branch Control: Take Branch=%0b, Target Address=0x%0h, Branch Type=%0b, PC+4=0x%h", 
                  dut.id_take_branch,
                  dut.id_branch_target_addr,
                  dut.id_stage_inst.branch_type,
                  dut.id_next_pc);         

        $display("EX: ALUSrcA=%0b, ALUinputA=%0d, ALUinputB=%0d, Shamt=0x%h, ALUControl=%0d, ALUResult=%0d, RD=%0d, RegWrite=%0b",
                 dut.ex_stage_inst.i_alu_src_a,
                 dut.ex_stage_inst.alu_input_a,
                 dut.ex_stage_inst.alu_input_b, 
                 dut.ex_stage_inst.i_shamt,
                 dut.ex_stage_inst.alu_control,
                 dut.ex_alu_result,
                 dut.ex_write_register,
                 dut.ex_reg_write);
        
        // Mostrar también los registros de origen y destino relevantes
        $display("REGS: Rs=%0d, Rt=%0d, MEM_Rd=%0d, WB_Rd=%0d", 
                 dut.ex_rs,
                 dut.ex_rt,
                 dut.mem_write_register,
                 dut.wb_write_register_out);
               
        $display("MEM: ALUResult=%0d, MemWrite=%0b, MemRead=%0b, RegWrite=%0b", 
                 dut.mem_alu_result,
                 dut.mem_mem_write,
                 dut.mem_mem_read,
                 dut.mem_reg_write_out);
                 
        $display("WB: WriteReg=%0d, WriteData=%0d, RegWrite=%0b", 
                 dut.wb_write_register_out,
                 dut.wb_write_data,
                 dut.wb_reg_write_out);
    end
  end
  
  // Ya no necesitamos la verificación basada en ciclos, 
  // ya que ahora se ejecuta cuando halt=1

  // Para generar formas de onda (VCD)
  initial begin
    $dumpfile("mips_simple.vcd");
    $dumpvars(0, mips_simple_tb);
  end

endmodule
